library verilog;
use verilog.vl_types.all;
entity bit_counter_vlg_vec_tst is
end bit_counter_vlg_vec_tst;
