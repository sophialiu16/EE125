library verilog;
use verilog.vl_types.all;
entity synch_counter_vlg_vec_tst is
end synch_counter_vlg_vec_tst;
