library verilog;
use verilog.vl_types.all;
entity abs_difference_calculator_vlg_vec_tst is
end abs_difference_calculator_vlg_vec_tst;
