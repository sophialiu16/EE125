library verilog;
use verilog.vl_types.all;
entity synch_counter_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end synch_counter_vlg_sample_tst;
