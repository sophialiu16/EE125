library verilog;
use verilog.vl_types.all;
entity guess_the_circuit_vlg_check_tst is
    port(
        y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end guess_the_circuit_vlg_check_tst;
