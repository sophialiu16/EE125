library verilog;
use verilog.vl_types.all;
entity kitchen_ctr_vlg_vec_tst is
end kitchen_ctr_vlg_vec_tst;
