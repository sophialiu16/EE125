library verilog;
use verilog.vl_types.all;
entity test_nat_therm_vlg_vec_tst is
end test_nat_therm_vlg_vec_tst;
