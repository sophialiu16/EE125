library verilog;
use verilog.vl_types.all;
entity guess_the_circuit_vlg_vec_tst is
end guess_the_circuit_vlg_vec_tst;
