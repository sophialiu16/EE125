library verilog;
use verilog.vl_types.all;
entity guess_the_circuit_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end guess_the_circuit_vlg_sample_tst;
