library verilog;
use verilog.vl_types.all;
entity calc_ceil_log2_vlg_vec_tst is
end calc_ceil_log2_vlg_vec_tst;
